LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Lab2Parte1 IS
PORT( 
SW : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END Lab2Parte1;

ARCHITECTURE Behavior OF Lab2Parte1 IS
BEGIN

HEX0 <= "1000000" WHEN SW = "00000" OR SW = "01010" OR SW = "10100" OR SW = "11110" ELSE
			"1111001" WHEN SW = "00001" OR SW = "01011" OR SW = "10101" OR SW = "11111" ELSE
			"0100100" WHEN SW = "00010" OR SW = "01100" OR SW = "10110" ELSE
			"0110000" WHEN SW = "00011" OR SW = "01101" OR SW = "10111" ELSE
			"0011001" WHEN SW = "00100" OR SW = "01110" OR SW = "11000" ELSE
			"0010010" WHEN SW = "00101" OR SW = "01111" OR SW = "11001" ELSE
			"0000010" WHEN SW = "00110" OR SW = "10000" OR SW = "11010" ELSE
			"1111000" WHEN SW = "00111" OR SW = "10001" OR SW = "11011" ELSE
			"0000000" WHEN SW = "01000" OR SW = "10010" OR SW = "11100" ELSE
			"0010000" WHEN SW = "01001" OR SW = "10011" OR SW = "11101" ELSE
			"1111111";
 
HEX1 <=   "0110000" WHEN SW >= "11110" ELSE
			 "0100100" WHEN SW >= "10100" ELSE
			 "1111001" WHEN SW >= "01010" ELSE
			 "1000000";
 
 
END Behavior;